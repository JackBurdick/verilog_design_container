module mux_4to1_df(Out, In, Sel)
output Out;
input [3:0]In;
input [1:0]Sel;